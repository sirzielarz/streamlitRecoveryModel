���      �sklearn.linear_model._logistic��LogisticRegression���)��}�(�penalty��l2��dual���tol�G?6��C-�C�G?�      �fit_intercept���intercept_scaling�K�class_weight�N�random_state�N�solver��lbfgs��max_iter�Kd�multi_class��auto��verbose�K �
warm_start���n_jobs�N�l1_ratio�N�n_features_in_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�n_iter_�hhK ��h ��R�(KK��h%�i4�����R�(Kh)NNNJ����J����K t�b�C8   �t�b�coef_�hhK ��h ��R�(KKK��h%�f8�����R�(Kh)NNNJ����J����K t�b�C D�i�@F�n͙k?��aq-��?���k0���t�b�
intercept_�hhK ��h ��R�(KK��h?�C��4=�濔t�b�_sklearn_version��0.24.1�ub.